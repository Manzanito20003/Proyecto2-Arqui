module hazard();
  
endmodule